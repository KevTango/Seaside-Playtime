library IEEE;
use  IEEE.STD_LOGIC_1164.all;
use  IEEE.STD_LOGIC_ARITH.all;
use  IEEE.STD_LOGIC_UNSIGNED.all;

entity score_disp_selector is
	port(
		Clk  : in std_logic;
		Ones : in std_logic_vector(5 downto 0);
		Tens : in std_logic_vector(5 downto 0);
		Hundreds : in std_logic_vector(5 downto 0);
		Thousands : in std_logic_vector(5 downto 0);
		pixel_row, pixel_column : in std_logic_vector (10 downto 0);
		score_output : out std_logic_vector(5 downto 0);
		score_enable : out std_logic
	);
end entity score_disp_selector;

architecture behaviour of score_disp_selector is
begin
	process(Clk, pixel_row, pixel_column, thousands, hundreds, tens, ones)
	begin 
		if (pixel_row >= 16 and pixel_row < 32 and pixel_column > 0 and pixel_column < 16) then
			score_output <= thousands;
			score_enable <= '1';
		elsif (pixel_row >= 16 and pixel_row < 32 and pixel_column >= 16 and pixel_column < 32) then
			score_output <= hundreds;
			score_enable <= '1';
		elsif (pixel_row >= 16 and pixel_row < 32 and pixel_column >= 32 and pixel_column < 48) then
			score_output <= tens;
			score_enable <= '1';
		elsif (pixel_row >= 16 and pixel_row < 32 and pixel_column >= 48 and pixel_column < 64) then
			score_output <= ones;
			score_enable <= '1';
		else
			score_output <= "000000";
			score_enable <= '0';
		end if;
	end process;
end architecture behaviour;
		